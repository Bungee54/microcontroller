-- Evan Allen, 9/7/2018

library IEEE;
use IEEE.numeric_std.all;

package microcontroller_package is
    constant word_size : NATURAL := 16;
    constant addr_size : NATURAL := word_size;
end microcontroller_package;